`include "define.vh"

module top (

// LEDs
output [3:0]    LED,

// USB3 FT601 Interface
input           ftdi_clk,
input           ftdi_rxf_n,
input           ftdi_txe_n,
output          ftdi_oe_n,
output          ftdi_rd_n,
output          ftdi_wr_n,
input  [31:0]   ftdi_data_IN,
output [31:0]   ftdi_data_OUT,
output [31:0]   ftdi_data_OE,
input  [3:0]    ftdi_be_IN,
output [3:0]    ftdi_be_OUT,
output [3:0]    ftdi_be_OE,

// 100MHz clock for USB processing
input           clk_100,

// DDR Interface
input           axi0_ACLK,
output          axi0_ARESETn,
output          axi0_ARQOS,
output          axi0_AWQOS,
output [5:0]    axi0_AWID,
output [32:0]   axi0_AWADDR,
output [7:0]    axi0_AWLEN,
output [2:0]    axi0_AWSIZE,
output [1:0]    axi0_AWBURST,
output          axi0_AWVALID,
output [3:0]    axi0_AWCACHE,
output          axi0_AWCOBUF,
output          axi0_AWLOCK,
output          axi0_AWAPCMD,
output          axi0_AWALLSTRB,
output [5:0]    axi0_ARID,
output [32:0]   axi0_ARADDR,
output [7:0]    axi0_ARLEN,
output [2:0]    axi0_ARSIZE,
output [1:0]    axi0_ARBURST,
output          axi0_ARVALID,
output          axi0_ARLOCK,
output          axi0_ARAPCMD,
output          axi0_WLAST,
output          axi0_WVALID,
output [511:0]  axi0_WDATA,
output [63:0]   axi0_WSTRB,
output          axi0_BREADY,
output          axi0_RREADY,
input           axi0_AWREADY,
input           axi0_ARREADY,
input           axi0_WREADY,
input [5:0]     axi0_BID,
input [1:0]     axi0_BRESP,
input           axi0_BVALID,
input [5:0]     axi0_RID,
input           axi0_RLAST,
input           axi0_RVALID,
input [511:0]   axi0_RDATA,
input [1:0]     axi0_RRESP,

input           axi1_ACLK,
output          axi1_ARESETn,
output          axi1_ARQOS,
output          axi1_AWQOS,
output [5:0]    axi1_AWID,
output [32:0]   axi1_AWADDR,
output [7:0]    axi1_AWLEN,
output [2:0]    axi1_AWSIZE,
output [1:0]    axi1_AWBURST,
output          axi1_AWVALID,
output [3:0]    axi1_AWCACHE,
output          axi1_AWCOBUF,
output          axi1_AWLOCK,
output          axi1_AWAPCMD,
output          axi1_AWALLSTRB,
output [5:0]    axi1_ARID,
output [32:0]   axi1_ARADDR,
output [7:0]    axi1_ARLEN,
output [2:0]    axi1_ARSIZE,
output [1:0]    axi1_ARBURST,
output          axi1_ARVALID,
output          axi1_ARLOCK,
output          axi1_ARAPCMD,
output          axi1_WLAST,
output          axi1_WVALID,
output [511:0]  axi1_WDATA,
output [63:0]   axi1_WSTRB,
output          axi1_BREADY,
output          axi1_RREADY,
input           axi1_AWREADY,
input           axi1_ARREADY,
input           axi1_WREADY,
input [5:0]     axi1_BID,
input [1:0]     axi1_BRESP,
input           axi1_BVALID,
input [5:0]     axi1_RID,
input           axi1_RLAST,
input           axi1_RVALID,
input [511:0]   axi1_RDATA,
input [1:0]     axi1_RRESP,

output          cfg_sel,
output          cfg_start,
output          cfg_reset,
input           cfg_done,
output          phy_rstn,
output          ctrl_rstn,
input           ddr_pll_lock,
output          ddr_pll_rstn,
//config
input           regACLK,
output [14:0]   regARADDR,
output [5:0]    regARID,
output [7:0]    regARLEN,
output [2:0]    regARSIZE,
output [1:0]    regARBURST,
output          regARVALID,
input           regARREADY,
input [31:0]    regRDATA,
input           regRVALID,
input           regRLAST,
input [1:0]     regRRESP,
input [5:0]     regRID,
output          regRREADY,
output [14:0]   regAWADDR,
output [5:0]    regAWID,
output [7:0]    regAWLEN,
output [2:0]    regAWSIZE,
output [1:0]    regAWBURST,
output          regAWVALID,
input           regAWREADY,

output [31:0]   regWDATA,
output [3:0]    regWSTRB,
output          regWLAST,
output          regWVALID,
input           regWREADY,

output          regBREADY,
input [5:0]     regBID,
input [1:0]     regBRESP,
input           regBVALID,

output          regARESETn,

input           jtag_inst1_CAPTURE,
input           jtag_inst1_DRCK,
input           jtag_inst1_RESET,
input           jtag_inst1_RUNTEST,
input           jtag_inst1_SEL,
input           jtag_inst1_SHIFT,
input           jtag_inst1_TCK,
input           jtag_inst1_TDI,
input           jtag_inst1_TMS,
input           jtag_inst1_UPDATE,
output          jtag_inst1_TDO
);


tools_core core0(

// LEDs
.LED(LED),

// USB3 Interface
.ftdi_clk(ftdi_clk),
.ftdi_rxf_n(ftdi_rxf_n),
.ftdi_txe_n(ftdi_txe_n),
.ftdi_oe_n(ftdi_oe_n),
.ftdi_rd_n(ftdi_rd_n),
.ftdi_wr_n(ftdi_wr_n),
.ftdi_data_IN(ftdi_data_IN),
.ftdi_data_OUT(ftdi_data_OUT),
.ftdi_data_OE(ftdi_data_OE),
.ftdi_be_IN(ftdi_be_IN),
.ftdi_be_OUT(ftdi_be_OUT),
.ftdi_be_OE(ftdi_be_OE),

// DDR Interface
.axi0_ACLK(axi0_ACLK),
.axi0_ARESETn(axi0_ARESETn),
.axi0_ARQOS(axi0_ARQOS),
.axi0_AWQOS(axi0_AWQOS),
.axi0_AWID(axi0_AWID),
.axi0_AWADDR(axi0_AWADDR),
.axi0_AWLEN(axi0_AWLEN),
.axi0_AWSIZE(axi0_AWSIZE),
.axi0_AWBURST(axi0_AWBURST),
.axi0_AWVALID(axi0_AWVALID),
.axi0_AWCACHE(axi0_AWCACHE),
.axi0_AWCOBUF(axi0_AWCOBUF),
.axi0_AWLOCK(axi0_AWLOCK),
.axi0_AWAPCMD(axi0_AWAPCMD),
.axi0_AWALLSTRB(axi0_AWALLSTRB),
.axi0_ARID(axi0_ARID),
.axi0_ARADDR(axi0_ARADDR),
.axi0_ARLEN(axi0_ARLEN),
.axi0_ARSIZE(axi0_ARSIZE),
.axi0_ARBURST(axi0_ARBURST),
.axi0_ARVALID(axi0_ARVALID),
.axi0_ARLOCK(axi0_ARLOCK),
.axi0_ARAPCMD(axi0_ARAPCMD),
.axi0_WLAST(axi0_WLAST),
.axi0_WVALID(axi0_WVALID),
.axi0_WDATA(axi0_WDATA),
.axi0_WSTRB(axi0_WSTRB),
.axi0_BREADY(axi0_BREADY),
.axi0_RREADY(axi0_RREADY),
.axi0_AWREADY(axi0_AWREADY),
.axi0_ARREADY(axi0_ARREADY),
.axi0_WREADY(axi0_WREADY),
.axi0_BID(axi0_BID),
.axi0_BRESP(axi0_BRESP),
.axi0_BVALID(axi0_BVALID),
.axi0_RID(axi0_RID),
.axi0_RLAST(axi0_RLAST),
.axi0_RVALID(axi0_RVALID),
.axi0_RDATA(axi0_RDATA),
.axi0_RRESP(axi0_RRESP),

.axi1_ACLK(axi1_ACLK),
.axi1_ARESETn(axi1_ARESETn),
.axi1_ARQOS(axi1_ARQOS),
.axi1_AWQOS(axi1_AWQOS),
.axi1_AWID(axi1_AWID),
.axi1_AWADDR(axi1_AWADDR),
.axi1_AWLEN(axi1_AWLEN),
.axi1_AWSIZE(axi1_AWSIZE),
.axi1_AWBURST(axi1_AWBURST),
.axi1_AWVALID(axi1_AWVALID),
.axi1_AWCACHE(axi1_AWCACHE),
.axi1_AWCOBUF(axi1_AWCOBUF),
.axi1_AWLOCK(axi1_AWLOCK),
.axi1_AWAPCMD(axi1_AWAPCMD),
.axi1_AWALLSTRB(axi1_AWALLSTRB),
.axi1_ARID(axi1_ARID),
.axi1_ARADDR(axi1_ARADDR),
.axi1_ARLEN(axi1_ARLEN),
.axi1_ARSIZE(axi1_ARSIZE),
.axi1_ARBURST(axi1_ARBURST),
.axi1_ARVALID(axi1_ARVALID),
.axi1_ARLOCK(axi1_ARLOCK),
.axi1_ARAPCMD(axi1_ARAPCMD),
.axi1_WLAST(axi1_WLAST),
.axi1_WVALID(axi1_WVALID),
.axi1_WDATA(axi1_WDATA),
.axi1_WSTRB(axi1_WSTRB),
.axi1_BREADY(axi1_BREADY),
.axi1_RREADY(axi1_RREADY),
.axi1_AWREADY(axi1_AWREADY),
.axi1_ARREADY(axi1_ARREADY),
.axi1_WREADY(axi1_WREADY),
.axi1_BID(axi1_BID),
.axi1_BRESP(axi1_BRESP),
.axi1_BVALID(axi1_BVALID),
.axi1_RID(axi1_RID),
.axi1_RLAST(axi1_RLAST),
.axi1_RVALID(axi1_RVALID),
.axi1_RDATA(axi1_RDATA),
.axi1_RRESP(axi1_RRESP),

.cfg_sel(cfg_sel),
.cfg_start(cfg_start),
.cfg_reset(cfg_reset),
.cfg_done(cfg_done),
.phy_rstn(phy_rstn),
.ctrl_rstn(ctrl_rstn),
.ddr_pll_lock(ddr_pll_lock),
.ddr_pll_rstn(ddr_pll_rstn),

.regACLK(regACLK),
.regARADDR(regARADDR),
.regARID(regARID),
.regARLEN(regARLEN),
.regARSIZE(regARSIZE),
.regARBURST(regARBURST),
.regARVALID(regARVALID),
.regARREADY(regARREADY),
.regRDATA(regRDATA),
.regRVALID(regRVALID),
.regRLAST(regRLAST),
.regRRESP(regRRESP),
.regRID(regRID),
.regRREADY(regRREADY),
.regAWADDR(regAWADDR),
.regAWID(regAWID),
.regAWLEN(regAWLEN),
.regAWSIZE(regAWSIZE),
.regAWBURST(regAWBURST),
.regAWVALID(regAWVALID),
.regAWREADY(regAWREADY),

.regWDATA(regWDATA),
.regWSTRB(regWSTRB),
.regWLAST(regWLAST),
.regWVALID(regWVALID),
.regWREADY(regWREADY),

.regBREADY(regBREADY),
.regBID(regBID),
.regBRESP(regBRESP),
.regBVALID(regBVALID),

.regARESETn(regARESETn),

.jtag_inst1_CAPTURE(jtag_inst1_CAPTURE),
.jtag_inst1_DRCK(jtag_inst1_DRCK),
.jtag_inst1_RESET(jtag_inst1_RESET),
.jtag_inst1_RUNTEST(jtag_inst1_RUNTEST),
.jtag_inst1_SEL(jtag_inst1_SEL),
.jtag_inst1_SHIFT(jtag_inst1_SHIFT),
.jtag_inst1_TCK(jtag_inst1_TCK),
.jtag_inst1_TDI(jtag_inst1_TDI),
.jtag_inst1_TMS(jtag_inst1_TMS),
.jtag_inst1_UPDATE(jtag_inst1_UPDATE),
.jtag_inst1_TDO(jtag_inst1_TDO)
);

endmodule