`define DBG_ID_WIDTH 4
`define CS_WIDTH (1<<`DBG_ID_WIDTH)-1
`define DR_WIDTH  82