
// Efinity Top-level template
// Version: 2025.1.110.5.9
// Date: 2025-11-12 23:50

// Copyright (C) 2013 - 2025 Efinix Inc. All rights reserved.

// This file may be used as a starting point for Efinity synthesis top-level target.
// The port list here matches what is expected by Efinity constraint files generated
// by the Efinity Interface Designer.

// To use this:
//     #1)  Save this file with a different name to a different directory, where source files are kept.
//              Example: you may wish to save as tools_core.v
//     #2)  Add the newly saved file into Efinity project as design file
//     #3)  Edit the top level entity in Efinity project to:  tools_core
//     #4)  Insert design content.


module tools_core
(
  (* syn_peri_port = 0 *) input ddr_pllin,
  (* syn_peri_port = 0 *) input ddr_pll_lock,
  (* syn_peri_port = 0 *) input regACLK,
  (* syn_peri_port = 0 *) input axi1_ACLK,
  (* syn_peri_port = 0 *) input axi0_ACLK,
  (* syn_peri_port = 0 *) input jtag_inst1_CAPTURE,
  (* syn_peri_port = 0 *) input jtag_inst1_DRCK,
  (* syn_peri_port = 0 *) input jtag_inst1_RESET,
  (* syn_peri_port = 0 *) input jtag_inst1_RUNTEST,
  (* syn_peri_port = 0 *) input jtag_inst1_SEL,
  (* syn_peri_port = 0 *) input jtag_inst1_SHIFT,
  (* syn_peri_port = 0 *) input jtag_inst1_TCK,
  (* syn_peri_port = 0 *) input jtag_inst1_TDI,
  (* syn_peri_port = 0 *) input jtag_inst1_TMS,
  (* syn_peri_port = 0 *) input jtag_inst1_UPDATE,
  (* syn_peri_port = 0 *) input axi0_ARREADY,
  (* syn_peri_port = 0 *) input axi1_ARREADY,
  (* syn_peri_port = 0 *) input axi0_AWREADY,
  (* syn_peri_port = 0 *) input axi1_AWREADY,
  (* syn_peri_port = 0 *) input [5:0] axi0_BID,
  (* syn_peri_port = 0 *) input [5:0] axi1_BID,
  (* syn_peri_port = 0 *) input [1:0] axi0_BRESP,
  (* syn_peri_port = 0 *) input [1:0] axi1_BRESP,
  (* syn_peri_port = 0 *) input axi0_BVALID,
  (* syn_peri_port = 0 *) input axi1_BVALID,
  (* syn_peri_port = 0 *) input cfg_done,
  (* syn_peri_port = 0 *) input regARREADY,
  (* syn_peri_port = 0 *) input regAWREADY,
  (* syn_peri_port = 0 *) input [5:0] regBID,
  (* syn_peri_port = 0 *) input [1:0] regBRESP,
  (* syn_peri_port = 0 *) input regBVALID,
  (* syn_peri_port = 0 *) input [31:0] regRDATA,
  (* syn_peri_port = 0 *) input [5:0] regRID,
  (* syn_peri_port = 0 *) input regRLAST,
  (* syn_peri_port = 0 *) input [1:0] regRRESP,
  (* syn_peri_port = 0 *) input regRVALID,
  (* syn_peri_port = 0 *) input regWREADY,
  (* syn_peri_port = 0 *) input [511:0] axi0_RDATA,
  (* syn_peri_port = 0 *) input [511:0] axi1_RDATA,
  (* syn_peri_port = 0 *) input [5:0] axi0_RID,
  (* syn_peri_port = 0 *) input [5:0] axi1_RID,
  (* syn_peri_port = 0 *) input axi0_RLAST,
  (* syn_peri_port = 0 *) input axi1_RLAST,
  (* syn_peri_port = 0 *) input [1:0] axi0_RRESP,
  (* syn_peri_port = 0 *) input [1:0] axi1_RRESP,
  (* syn_peri_port = 0 *) input axi0_RVALID,
  (* syn_peri_port = 0 *) input axi1_RVALID,
  (* syn_peri_port = 0 *) input axi0_WREADY,
  (* syn_peri_port = 0 *) input axi1_WREADY,
  (* syn_peri_port = 0 *) output ddr_pll_rstn,
  (* syn_peri_port = 0 *) output jtag_inst1_TDO,
  (* syn_peri_port = 0 *) output [32:0] axi0_ARADDR,
  (* syn_peri_port = 0 *) output [32:0] axi1_ARADDR,
  (* syn_peri_port = 0 *) output axi0_ARAPCMD,
  (* syn_peri_port = 0 *) output axi1_ARAPCMD,
  (* syn_peri_port = 0 *) output [1:0] axi0_ARBURST,
  (* syn_peri_port = 0 *) output [1:0] axi1_ARBURST,
  (* syn_peri_port = 0 *) output [5:0] axi0_ARID,
  (* syn_peri_port = 0 *) output [5:0] axi1_ARID,
  (* syn_peri_port = 0 *) output [7:0] axi0_ARLEN,
  (* syn_peri_port = 0 *) output [7:0] axi1_ARLEN,
  (* syn_peri_port = 0 *) output axi0_ARLOCK,
  (* syn_peri_port = 0 *) output axi1_ARLOCK,
  (* syn_peri_port = 0 *) output axi0_ARQOS,
  (* syn_peri_port = 0 *) output axi1_ARQOS,
  (* syn_peri_port = 0 *) output [2:0] axi0_ARSIZE,
  (* syn_peri_port = 0 *) output [2:0] axi1_ARSIZE,
  (* syn_peri_port = 0 *) output axi0_ARESETn,
  (* syn_peri_port = 0 *) output axi1_ARESETn,
  (* syn_peri_port = 0 *) output axi0_ARVALID,
  (* syn_peri_port = 0 *) output axi1_ARVALID,
  (* syn_peri_port = 0 *) output [32:0] axi0_AWADDR,
  (* syn_peri_port = 0 *) output [32:0] axi1_AWADDR,
  (* syn_peri_port = 0 *) output axi0_AWALLSTRB,
  (* syn_peri_port = 0 *) output axi1_AWALLSTRB,
  (* syn_peri_port = 0 *) output axi0_AWAPCMD,
  (* syn_peri_port = 0 *) output axi1_AWAPCMD,
  (* syn_peri_port = 0 *) output [1:0] axi0_AWBURST,
  (* syn_peri_port = 0 *) output [1:0] axi1_AWBURST,
  (* syn_peri_port = 0 *) output [3:0] axi0_AWCACHE,
  (* syn_peri_port = 0 *) output [3:0] axi1_AWCACHE,
  (* syn_peri_port = 0 *) output axi0_AWCOBUF,
  (* syn_peri_port = 0 *) output axi1_AWCOBUF,
  (* syn_peri_port = 0 *) output [5:0] axi0_AWID,
  (* syn_peri_port = 0 *) output [5:0] axi1_AWID,
  (* syn_peri_port = 0 *) output [7:0] axi0_AWLEN,
  (* syn_peri_port = 0 *) output [7:0] axi1_AWLEN,
  (* syn_peri_port = 0 *) output axi0_AWLOCK,
  (* syn_peri_port = 0 *) output axi1_AWLOCK,
  (* syn_peri_port = 0 *) output axi0_AWQOS,
  (* syn_peri_port = 0 *) output axi1_AWQOS,
  (* syn_peri_port = 0 *) output [2:0] axi0_AWSIZE,
  (* syn_peri_port = 0 *) output [2:0] axi1_AWSIZE,
  (* syn_peri_port = 0 *) output axi0_AWVALID,
  (* syn_peri_port = 0 *) output axi1_AWVALID,
  (* syn_peri_port = 0 *) output axi0_BREADY,
  (* syn_peri_port = 0 *) output axi1_BREADY,
  (* syn_peri_port = 0 *) output phy_rstn,
  (* syn_peri_port = 0 *) output cfg_reset,
  (* syn_peri_port = 0 *) output cfg_sel,
  (* syn_peri_port = 0 *) output cfg_start,
  (* syn_peri_port = 0 *) output [14:0] regARADDR,
  (* syn_peri_port = 0 *) output [1:0] regARBURST,
  (* syn_peri_port = 0 *) output regARESETn,
  (* syn_peri_port = 0 *) output [5:0] regARID,
  (* syn_peri_port = 0 *) output [7:0] regARLEN,
  (* syn_peri_port = 0 *) output [2:0] regARSIZE,
  (* syn_peri_port = 0 *) output regARVALID,
  (* syn_peri_port = 0 *) output [14:0] regAWADDR,
  (* syn_peri_port = 0 *) output [1:0] regAWBURST,
  (* syn_peri_port = 0 *) output [5:0] regAWID,
  (* syn_peri_port = 0 *) output [7:0] regAWLEN,
  (* syn_peri_port = 0 *) output [2:0] regAWSIZE,
  (* syn_peri_port = 0 *) output regAWVALID,
  (* syn_peri_port = 0 *) output regBREADY,
  (* syn_peri_port = 0 *) output regRREADY,
  (* syn_peri_port = 0 *) output [31:0] regWDATA,
  (* syn_peri_port = 0 *) output regWLAST,
  (* syn_peri_port = 0 *) output [3:0] regWSTRB,
  (* syn_peri_port = 0 *) output regWVALID,
  (* syn_peri_port = 0 *) output ctrl_rstn,
  (* syn_peri_port = 0 *) output axi0_RREADY,
  (* syn_peri_port = 0 *) output axi1_RREADY,
  (* syn_peri_port = 0 *) output [511:0] axi0_WDATA,
  (* syn_peri_port = 0 *) output [511:0] axi1_WDATA,
  (* syn_peri_port = 0 *) output axi0_WLAST,
  (* syn_peri_port = 0 *) output axi1_WLAST,
  (* syn_peri_port = 0 *) output [63:0] axi0_WSTRB,
  (* syn_peri_port = 0 *) output [63:0] axi1_WSTRB,
  (* syn_peri_port = 0 *) output axi0_WVALID,
  (* syn_peri_port = 0 *) output axi1_WVALID
);


endmodule

